LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DFF IS PORT (
		D, Clock: IN STD_LOGIC;
		Q: OUT STD_LOGIC);
END DFF;

ARCHITECTURE Behavior OF DFF IS
BEGIN
	PROCESS(Clock)
	BEGIN
		IF (Clock'Event AND Clock = '1') THEN
			Q <= D;
		END IF;
	END PROCESS;
END Behavior;